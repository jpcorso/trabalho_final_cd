library verilog;
use verilog.vl_types.all;
entity contador_top_vlg_vec_tst is
end contador_top_vlg_vec_tst;
